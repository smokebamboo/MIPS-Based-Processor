----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:22:58 03/16/2025 
-- Design Name: 
-- Module Name:    Adder_32_bit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Adder_32_bit is
    Port( Input : in  STD_LOGIC_VECTOR (31 downto 0);
          Output : out  STD_LOGIC_VECTOR (31 downto 0));
end Adder_32_bit;

architecture Behavioral of Adder_32_bit is

begin

	Output <= Input + "00000000000000000000000000000100";
	
end Behavioral;

